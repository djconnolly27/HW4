//------------------------------------------------------------------------------
// Test harness validates hw4testbench by connecting it to various functional
// or broken register files, and verifying that it correctly identifies each
//------------------------------------------------------------------------------

`include "regfile.v"

module hw4testbenchharness();

  wire[31:0]	ReadData1;	// Data from first register read
  wire[31:0]	ReadData2;	// Data from second register read
  wire[31:0]	WriteData;	// Data to write to register
  wire[4:0]	ReadRegister1;	// Address of first register to read
  wire[4:0]	ReadRegister2;	// Address of second register to read
  wire[4:0]	WriteRegister;  // Address of register to write
  wire		RegWrite;	// Enable writing of register when High
  wire		Clk;		// Clock (Positive Edge Triggered)

  reg		begintest;	// Set High to begin testing register file
  wire  	endtest;    	// Set High to signal test completion
  wire		dutpassed;	// Indicates whether register file passed tests

  // Instantiate the register file being tested.  DUT = Device Under Test
  regfile DUT
  (
    .ReadData1(ReadData1),
    .ReadData2(ReadData2),
    .WriteData(WriteData),
    .ReadRegister1(ReadRegister1),
    .ReadRegister2(ReadRegister2),
    .WriteRegister(WriteRegister),
    .RegWrite(RegWrite),
    .Clk(Clk)
  );

  // Instantiate test bench to test the DUT
  hw4testbench tester
  (
    .begintest(begintest),
    .endtest(endtest),
    .dutpassed(dutpassed),
    .ReadData1(ReadData1),
    .ReadData2(ReadData2),
    .WriteData(WriteData),
    .ReadRegister1(ReadRegister1),
    .ReadRegister2(ReadRegister2),
    .WriteRegister(WriteRegister),
    .RegWrite(RegWrite),
    .Clk(Clk)
  );

  // Test harness asserts 'begintest' for 1000 time steps, starting at time 10
  initial begin
    begintest=0;
    #10;
    begintest=1;
    #1000;
  end

  // Display test results ('dutpassed' signal) once 'endtest' goes high
  always @(posedge endtest) begin
    $display("DUT passed?: %b", dutpassed);
  end

endmodule


//------------------------------------------------------------------------------
// Your HW4 test bench
//   Generates signals to drive register file and passes them back up one
//   layer to the test harness. This lets us plug in various working and
//   broken register files to test.
//
//   Once 'begintest' is asserted, begin testing the register file.
//   Once your test is conclusive, set 'dutpassed' appropriately and then
//   raise 'endtest'.
//------------------------------------------------------------------------------

module hw4testbench
(
// Test bench driver signal connections
input	   		begintest,	// Triggers start of testing
output reg 		endtest,	// Raise once test completes
output reg 		dutpassed,	// Signal test result

// Register File DUT connections
input[31:0]		ReadData1,
input[31:0]		ReadData2,
output reg[31:0]	WriteData,
output reg[4:0]		ReadRegister1,
output reg[4:0]		ReadRegister2,
output reg[4:0]		WriteRegister,
output reg		RegWrite,
output reg		Clk
);

  // Initialize register driver signals
  initial begin
    WriteData=32'd0;
    ReadRegister1=5'd0;
    ReadRegister2=5'd0;
    WriteRegister=5'd0;
    RegWrite=0;
    Clk=0;
  end

  integer address, index;

  task reset_registers;
    for(address = 0; address < 32; address = address + 1) begin
      WriteRegister=address;
      WriteData=32'd0;
      RegWrite=1;
      #5 Clk=1; #5 Clk=0; #5 Clk=1; #5 Clk=0;
    end
  endtask

  // Once 'begintest' is asserted, start running test cases
  always @(posedge begintest) begin
    endtest = 0;
    dutpassed = 1;
    #10

  // Test Case 1:
  //   Write '42' to register 2, verify with Read Ports 1 and 2
  reset_registers();
  WriteRegister = 5'd2;
  WriteData = 32'd42;
  RegWrite = 1;
  ReadRegister1 = 5'd2;
  ReadRegister2 = 5'd2;
  #5 Clk=1; #5 Clk=0;	// Generate single clock pulse

  // Verify expectations and report test result
  if((ReadData1 !== 42) || (ReadData2 !== 42)) begin
    dutpassed = 0;	// Set to 'false' on failure
    $display("Test Case 1 Failed");
  end

  // Test Case 2:
  //   Write '15' to register 2, verify with Read Ports 1 and 2
  reset_registers();
  WriteRegister = 5'd2;
  WriteData = 32'd15;
  RegWrite = 1;
  ReadRegister1 = 5'd2;
  ReadRegister2 = 5'd2;
  #5 Clk=1; #5 Clk=0;

  if((ReadData1 !== 15) || (ReadData2 !== 15)) begin
    dutpassed = 0;
    $display("Test Case 2 Failed");
  end


  // Test Case 3:
  //   Turn off write enable
  //   Write '11' to register a random register, verify that all registers were not written to with Read Ports 1 and 2
  reset_registers();
  WriteRegister = $random%31+1;
  WriteData = 32'd11;
  RegWrite = 0;
  for(index=0;index <=15;index = index + 1) begin
    ReadRegister1 = index;
    ReadRegister2 = index + 16;
    #5 Clk=1; #5 Clk=0;

    // The value in register 2 should not have changed from the last test, and should still read 15
    if((ReadData1 !== 0) || (ReadData2 !== 0)) begin
      dutpassed = 0;
      $display("Test Case 3 Failed");
    end
  end

  // Test Case 4:
  //   Turn on write enable
  //   Write '23' to register 0, verify that the register 0 still reads
  //    the constant value 0 with Read Ports 1 and 2
  reset_registers();
  WriteRegister = 5'd0;
  WriteData = 32'd23;
  RegWrite = 1;
  ReadRegister1 = 5'd0;
  ReadRegister2 = 5'd0;
  #5 Clk=1; #5 Clk=0;

  if((ReadData1 !== 0) || (ReadData2 !== 0)) begin
    dutpassed = 0;
    $display("Test Case 4 Failed");
  end

  // Test Case 5:
  //   Turn on write enable
  //   Write '23' to register 8, verify that register 8 reads '23'
  //    and that register 4 still reads zero. This verifies the decoder is working
  reset_registers();
  WriteRegister = 5'd8;
  WriteData = 32'd23;
  RegWrite = 1;
  ReadRegister1 = 5'd8;
  ReadRegister2 = 5'd4;
  #5 Clk=1; #5 Clk=0;

  if((ReadData1 !== 23) || (ReadData2 !== 0)) begin
    dutpassed = 0;
    $display("Test Case 5 Failed");
  end

  // Test Case 6:
  //   Turn on write enable
  //   Write '9' to register 6, verify that register 22 reads '0' and is unaffected
  //    and that register 31 reads '0' is unaffected
  reset_registers();
  WriteRegister = 5'd6;
  WriteData = 32'd9;
  RegWrite = 1;
  ReadRegister1 = 5'd22;
  ReadRegister2 = 5'd31;
  #5 Clk=1; #5 Clk=0;

  if((ReadData1 !== 0) || (ReadData2 !== 0)) begin
    dutpassed = 0;
    $display("Test Case 6 Failed");
  end

  // Test Case 7:
  //   Turn on write enable
  //   Checks that nothing is written until after a positive clock edge occurs
  reset_registers();
  WriteRegister = 5'd8;
  WriteData = 32'd9;
  RegWrite = 1;
  ReadRegister1 = 5'd8;
  ReadRegister2 = 5'd8;

  if((ReadData1 !== 0) || (ReadData2 !== 0)) begin
    dutpassed = 0;
    $display("Test Case 7, Part 1 Failed");
  end

  #5 Clk=1; #5 Clk=0;
  if((ReadData1 !== 9) || (ReadData2 !== 9)) begin
    dutpassed = 0;
    $display("Test Case 7, Part 2 Failed");
  end

  // Test Case 8:
  //   Write to a random port
  //   Check the values of all ports
  reset_registers();
  WriteRegister = $random%31+1;
  WriteData = 32'd9;
  RegWrite = 1;
  for(index=0;index <= 15;index = index + 1) begin
    ReadRegister1 = index+16;
    ReadRegister2 = index+16;
    #5 Clk=1; #5 Clk=0;

    if(((ReadRegister1 == WriteRegister) && (ReadData1 !== 9)) || ((ReadRegister2 == WriteRegister) && (ReadData2 !== 9)) || ((ReadRegister1 !== WriteRegister) && (ReadData1 !== 0)) || ((ReadRegister1 !== WriteRegister) && (ReadData1 !== 0))) begin
      dutpassed = 0;
      $display("Test Case 8 Failed");
    end
  end


  // All done!  Wait a moment and signal test completion.
  #5
  endtest = 1;

end

endmodule
